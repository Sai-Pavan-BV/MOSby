module pc();
endmodule