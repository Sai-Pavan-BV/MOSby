module inst_cache (
    ports
);
    
endmodule